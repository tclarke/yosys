(* techmap_celltype = "C" *)
module __C_0805_2012Metric #(
  parameter layer="F.Cu",
  parameter reference="REF**",
  parameter value="C_0805_2012Metric")
  (inout A, inout B);

  (* layer = layer *)
  (* reference = reference *)
  (* value = value *)
  (* footprint = "Capacitor_SMD:C_0805_2012Metric" *)
  C_0805_2012Metric __cell(A, B);


endmodule